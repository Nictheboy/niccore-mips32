/* 
 *  Description : Full 32-bit Carry-Lookahead Adder.
 *  Author      : nictheboy <nictheboy@outlook.com>
 *  Create Date : 2025/10/11 
 * 
 */

module adder (
    input  [31:0] a,
    input  [31:0] b,
    output [31:0] sum
);
    wire [31:0] c;
    assign c[0] = (a[0] & b[0]);
    assign c[1] = (a[1] & b[1]) | ((a[0] & b[0]) & (a[1] | b[1]));
    assign c[2] = (a[2] & b[2]) | ((a[1] & b[1]) & (a[2] | b[2])) | ((a[0] & b[0]) & (a[1] | b[1]) & (a[2] | b[2]));
    assign c[3] = (a[3] & b[3]) | ((a[2] & b[2]) & (a[3] | b[3])) | ((a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3])) | ((a[0] & b[0]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]));
    assign c[4] = (a[4] & b[4]) | ((a[3] & b[3]) & (a[4] | b[4])) | ((a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4])) | ((a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4])) | ((a[0] & b[0]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]));
    assign c[5] = (a[5] & b[5]) | ((a[4] & b[4]) & (a[5] | b[5])) | ((a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5])) | ((a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5])) | ((a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5])) | ((a[0] & b[0]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]));
    assign c[6] = (a[6] & b[6]) | ((a[5] & b[5]) & (a[6] | b[6])) | ((a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6])) | ((a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6])) | ((a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6])) | ((a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6])) | ((a[0] & b[0]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]));
    assign c[7] = (a[7] & b[7]) | ((a[6] & b[6]) & (a[7] | b[7])) | ((a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7])) | ((a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7])) | ((a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7])) | ((a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7])) | ((a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7])) | ((a[0] & b[0]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]));
    assign c[8] = (a[8] & b[8]) | ((a[7] & b[7]) & (a[8] | b[8])) | ((a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8])) | ((a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8])) | ((a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8])) | ((a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8])) | ((a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8])) | ((a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8])) | ((a[0] & b[0]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]));
    assign c[9] = (a[9] & b[9]) | ((a[8] & b[8]) & (a[9] | b[9])) | ((a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[10] = (a[10] & b[10]) | ((a[10] | b[10]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[11] = (a[11] & b[11]) | ((a[10] & b[10]) & (a[11] | b[11])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[12] = (a[12] & b[12]) | ((a[11] & b[11]) & (a[12] | b[12])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[13] = (a[13] & b[13]) | ((a[12] & b[12]) & (a[13] | b[13])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[14] = (a[14] & b[14]) | ((a[13] & b[13]) & (a[14] | b[14])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[15] = (a[15] & b[15]) | ((a[14] & b[14]) & (a[15] | b[15])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[16] = (a[16] & b[16]) | ((a[15] & b[15]) & (a[16] | b[16])) | ((a[14] & b[14]) & (a[15] | b[15]) & (a[16] | b[16])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[17] = (a[17] & b[17]) | ((a[16] & b[16]) & (a[17] | b[17])) | ((a[15] & b[15]) & (a[16] | b[16]) & (a[17] | b[17])) | ((a[14] & b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[18] = (a[18] & b[18]) | ((a[17] & b[17]) & (a[18] | b[18])) | ((a[16] & b[16]) & (a[17] | b[17]) & (a[18] | b[18])) | ((a[15] & b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18])) | ((a[14] & b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[19] = (a[19] & b[19]) | ((a[18] & b[18]) & (a[19] | b[19])) | ((a[17] & b[17]) & (a[18] | b[18]) & (a[19] | b[19])) | ((a[16] & b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19])) | ((a[15] & b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19])) | ((a[14] & b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] & b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] | b[1]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[20] = (a[20] & b[20]) | ((a[19] & b[19]) & (a[20] | b[20])) | ((a[18] & b[18]) & (a[19] | b[19]) & (a[20] | b[20])) | ((a[17] & b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20])) | ((a[16] & b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20])) | ((a[15] & b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20])) | ((a[14] & b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] & b[1]) & (a[20] | b[20]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] | b[1]) & (a[20] | b[20]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[21] = (a[21] & b[21]) | ((a[20] & b[20]) & (a[21] | b[21])) | ((a[19] & b[19]) & (a[20] | b[20]) & (a[21] | b[21])) | ((a[18] & b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21])) | ((a[17] & b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21])) | ((a[16] & b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21])) | ((a[15] & b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21])) | ((a[14] & b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] & b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] | b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[22] = (a[22] & b[22]) | ((a[21] & b[21]) & (a[22] | b[22])) | ((a[20] & b[20]) & (a[21] | b[21]) & (a[22] | b[22])) | ((a[19] & b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22])) | ((a[18] & b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22])) | ((a[17] & b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22])) | ((a[16] & b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22])) | ((a[15] & b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22])) | ((a[14] & b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] & b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] | b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[23] = (a[23] & b[23]) | ((a[22] & b[22]) & (a[23] | b[23])) | ((a[21] & b[21]) & (a[22] | b[22]) & (a[23] | b[23])) | ((a[20] & b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23])) | ((a[19] & b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23])) | ((a[18] & b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23])) | ((a[17] & b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23])) | ((a[16] & b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23])) | ((a[15] & b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23])) | ((a[14] & b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] & b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] | b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[24] = (a[24] & b[24]) | ((a[23] & b[23]) & (a[24] | b[24])) | ((a[22] & b[22]) & (a[23] | b[23]) & (a[24] | b[24])) | ((a[21] & b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24])) | ((a[20] & b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24])) | ((a[19] & b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24])) | ((a[18] & b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24])) | ((a[17] & b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24])) | ((a[16] & b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24])) | ((a[15] & b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24])) | ((a[14] & b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] & b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] | b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[25] = (a[25] & b[25]) | ((a[24] & b[24]) & (a[25] | b[25])) | ((a[23] & b[23]) & (a[24] | b[24]) & (a[25] | b[25])) | ((a[22] & b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25])) | ((a[21] & b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25])) | ((a[20] & b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25])) | ((a[19] & b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25])) | ((a[18] & b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25])) | ((a[17] & b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25])) | ((a[16] & b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25])) | ((a[15] & b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25])) | ((a[14] & b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] & b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] | b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[26] = (a[26] & b[26]) | ((a[25] & b[25]) & (a[26] | b[26])) | ((a[24] & b[24]) & (a[25] | b[25]) & (a[26] | b[26])) | ((a[23] & b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26])) | ((a[22] & b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26])) | ((a[21] & b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26])) | ((a[20] & b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26])) | ((a[19] & b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26])) | ((a[18] & b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26])) | ((a[17] & b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26])) | ((a[16] & b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26])) | ((a[15] & b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26])) | ((a[14] & b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] & b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] | b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[27] = (a[27] & b[27]) | ((a[26] & b[26]) & (a[27] | b[27])) | ((a[25] & b[25]) & (a[26] | b[26]) & (a[27] | b[27])) | ((a[24] & b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27])) | ((a[23] & b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27])) | ((a[22] & b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27])) | ((a[21] & b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27])) | ((a[20] & b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27])) | ((a[19] & b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27])) | ((a[18] & b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27])) | ((a[17] & b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27])) | ((a[16] & b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27])) | ((a[15] & b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27])) | ((a[14] & b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] & b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] | b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[28] = (a[28] & b[28]) | ((a[27] & b[27]) & (a[28] | b[28])) | ((a[26] & b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[25] & b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[24] & b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[23] & b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[22] & b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[21] & b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[20] & b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[19] & b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[18] & b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[17] & b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[16] & b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[15] & b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[14] & b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] & b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] | b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[29] = (a[29] & b[29]) | ((a[28] & b[28]) & (a[29] | b[29])) | ((a[27] & b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[26] & b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[25] & b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[24] & b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[23] & b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[22] & b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[21] & b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[20] & b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[19] & b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[18] & b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[17] & b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[16] & b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[15] & b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[14] & b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[2] & b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] & b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] | b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[2] | b[2]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[30] = (a[30] & b[30]) | ((a[29] & b[29]) & (a[30] | b[30])) | ((a[28] & b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[27] & b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[26] & b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[25] & b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[24] & b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[23] & b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[22] & b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[21] & b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[20] & b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[19] & b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[18] & b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[17] & b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[16] & b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[15] & b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[14] & b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[2] & b[2]) & (a[30] | b[30]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] & b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[2] | b[2]) & (a[30] | b[30]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] | b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[2] | b[2]) & (a[30] | b[30]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign c[31] = (a[31] & b[31]) | ((a[30] & b[30]) & (a[31] | b[31])) | ((a[29] & b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[28] & b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[27] & b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[26] & b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[25] & b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[24] & b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[23] & b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[22] & b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[21] & b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[20] & b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[19] & b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[18] & b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[17] & b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[16] & b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[15] & b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[14] & b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[13] & b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[12] & b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[11] & b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[10] & b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31]) & (a[9] & b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31]) & (a[8] & b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31]) & (a[7] & b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31]) & (a[6] & b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31]) & (a[5] & b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31]) & (a[4] & b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[30] | b[30]) & (a[31] | b[31]) & (a[3] & b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[2] & b[2]) & (a[30] | b[30]) & (a[31] | b[31]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] & b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[2] | b[2]) & (a[30] | b[30]) & (a[31] | b[31]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9])) | ((a[0] & b[0]) & (a[10] | b[10]) & (a[11] | b[11]) & (a[12] | b[12]) & (a[13] | b[13]) & (a[14] | b[14]) & (a[15] | b[15]) & (a[16] | b[16]) & (a[17] | b[17]) & (a[18] | b[18]) & (a[19] | b[19]) & (a[1] | b[1]) & (a[20] | b[20]) & (a[21] | b[21]) & (a[22] | b[22]) & (a[23] | b[23]) & (a[24] | b[24]) & (a[25] | b[25]) & (a[26] | b[26]) & (a[27] | b[27]) & (a[28] | b[28]) & (a[29] | b[29]) & (a[2] | b[2]) & (a[30] | b[30]) & (a[31] | b[31]) & (a[3] | b[3]) & (a[4] | b[4]) & (a[5] | b[5]) & (a[6] | b[6]) & (a[7] | b[7]) & (a[8] | b[8]) & (a[9] | b[9]));
    assign sum = a ^ b ^ {c, 1'b0};
endmodule
